`timescale 1ns/1ps

module tb_can_error_handling;

  // DUT inputs
  logic clk;
  logic rst;
  logic rx_bit;
  logic tx_bit;
  logic tx_active;
  logic sample_point;
  logic bit_de_stuffing_ff;
  logic remove_stuff_bit;
  logic rx_bit_curr;
  logic rx_bit_prev;
  logic in_arbitration;
  logic in_ack_slot;
  logic in_crc_delimiter;
  logic in_ack_delimiter;
  logic in_eof;
  logic crc_check_done;
  logic crc_rx_valid;
  logic crc_rx_match;
  logic overload_request;
  logic dominant_after_flag;

  // DUT outputs
  logic bit_error;
  logic stuff_error;
  logic crc_error;
  logic form_error;
  logic ack_error;
  logic [7:0] tec;
  logic [7:0] rec;
  logic error_active;
  logic error_passive;
  logic bus_off;

  // Clock gen
  always #5 clk = ~clk;

  // DUT instance
  can_error_detection dut (
    .clk(clk),
    .rst(rst),
    .rx_bit(rx_bit),
    .tx_bit(tx_bit),
    .tx_active(tx_active),
    .sample_point(sample_point),
    .bit_de_stuffing_ff(bit_de_stuffing_ff),
    .remove_stuff_bit(remove_stuff_bit),
    .rx_bit_curr(rx_bit_curr),
    .rx_bit_prev(rx_bit_prev),
    .in_arbitration(in_arbitration),
    .in_ack_slot(in_ack_slot),
    .in_crc_delimiter(in_crc_delimiter),
    .in_ack_delimiter(in_ack_delimiter),
    .in_eof(in_eof),
    .crc_check_done(crc_check_done),
    .crc_rx_valid(crc_rx_valid),
    .crc_rx_match(crc_rx_match),
    .overload_request(overload_request),
    .dominant_after_flag(dominant_after_flag),
    .bit_error(bit_error),
    .stuff_error(stuff_error),
    .crc_error(crc_error),
    .form_error(form_error),
    .ack_error(ack_error),
    .tec(tec),
    .rec(rec),
    .error_active(error_active),
    .error_passive(error_passive),
    .bus_off(bus_off)
  );

  // Stimulus
  initial begin
    $monitor($time,,
      " rx=%0b tx=%0b bit_err=%0b stuff_err=%0b crc_err=%0b form_err=%0b ack_err=%0b tec=%0d rec=%0d act=%0b pas=%0b bus_off=%0b",
      rx_bit, tx_bit, bit_error, stuff_error, crc_error, form_error, ack_error,
      tec, rec, error_active, error_passive, bus_off);

    // Reset
    clk = 0;
    rst = 0;
    rx_bit = 1;
    tx_bit = 1;
    tx_active = 0;
    sample_point = 0;
    bit_de_stuffing_ff = 0;
    remove_stuff_bit   = 0;
    rx_bit_curr = 1;
    rx_bit_prev = 1;
    in_arbitration = 0;
    in_ack_slot = 0;
    in_crc_delimiter = 0;
    in_ack_delimiter = 0;
    in_eof = 0;
    crc_check_done = 0;
    crc_rx_valid = 0;
    crc_rx_match = 1;
    overload_request = 0;
    dominant_after_flag = 0;

    #20 rst = 1;

    // --- Trigger Bit Error ---
    #10 sample_point = 1;
        tx_active = 1;
        tx_bit = 1; rx_bit = 0;   // mismatch → bit_error
    #10 sample_point = 0; tx_active=0;

    // --- Trigger Stuff Error ---
    #20 sample_point = 1;
        bit_de_stuffing_ff = 1;
        remove_stuff_bit   = 1;
        rx_bit_curr = 0; rx_bit_prev = 0;
    #10 sample_point = 0;
        bit_de_stuffing_ff = 0; remove_stuff_bit = 0;

    // --- Trigger CRC Error ---
    #20 crc_check_done = 1; crc_rx_valid = 1; crc_rx_match = 0;
    #10 crc_check_done = 0;

    // --- Trigger Form Error ---
    #20 sample_point = 1; in_crc_delimiter = 1; rx_bit = 0;
    #10 sample_point = 0; in_crc_delimiter = 0; rx_bit = 1;

    // --- Trigger ACK Error ---
    #20 sample_point = 1; tx_active = 1; in_ack_slot = 1; rx_bit = 1;
    #10 sample_point = 0; in_ack_slot = 0;

    // Let counters update
    #100;

    $finish;
  end

endmodule
